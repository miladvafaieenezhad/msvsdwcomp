* SPICE3 file created from MY_INVERTER_0.ext - technology: sky130A

.subckt inverter_post_layout A VP Y VN

X0 Y A VN VN sky130_fd_pr__nfet_01v8  w=8.4 l=0.15

X1 VN A Y VN sky130_fd_pr__nfet_01v8  w=8.4 l=0.15

X2 Y A VP VP sky130_fd_pr__pfet_01v8 w=8.4 l=0.15

X3 VP A Y VP sky130_fd_pr__pfet_01v8 w=8.4 l=0.15

.ends
