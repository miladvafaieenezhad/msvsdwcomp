MACRO MY_RO
  ORIGIN 0 0 ;
  FOREIGN MY_RO 0 0 ;
  SIZE 5.16 BY 30.24 ;
  PIN VN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
      LAYER M3 ;
        RECT 1.58 3.595 1.86 3.965 ;
      LAYER M2 ;
        RECT 1.72 3.64 3.44 3.92 ;
      LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
      LAYER M3 ;
        RECT 2.87 15.8 3.15 22 ;
      LAYER M3 ;
        RECT 3.3 6.72 3.58 7.56 ;
      LAYER M2 ;
        RECT 3.01 7.42 3.44 7.7 ;
      LAYER M3 ;
        RECT 2.87 7.56 3.15 15.96 ;
    END
  END VN
  PIN VP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M3 ;
        RECT 1.58 11.155 1.86 11.525 ;
      LAYER M2 ;
        RECT 1.72 11.2 3.44 11.48 ;
      LAYER M3 ;
        RECT 3.3 11.155 3.58 11.525 ;
      LAYER M3 ;
        RECT 2.87 23.36 3.15 29.56 ;
      LAYER M3 ;
        RECT 1.58 14.28 1.86 22.68 ;
      LAYER M2 ;
        RECT 1.72 22.54 3.01 22.82 ;
      LAYER M3 ;
        RECT 2.87 22.68 3.15 23.52 ;
    END
  END VP
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
      LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
      LAYER M2 ;
        RECT 4.14 2.8 4.46 3.08 ;
      LAYER M3 ;
        RECT 4.16 2.94 4.44 12.18 ;
      LAYER M2 ;
        RECT 4.14 12.04 4.46 12.32 ;
    END
  END A
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.55 22.12 2.75 22.4 ;
      LAYER M2 ;
        RECT 1.55 22.96 2.75 23.24 ;
      LAYER M2 ;
        RECT 1.99 22.12 2.31 22.4 ;
      LAYER M3 ;
        RECT 2.01 22.26 2.29 23.1 ;
      LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
    END
  END Y
  OBS 
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.7 7 1.02 7.28 ;
  LAYER M3 ;
        RECT 0.72 7.14 1 7.98 ;
  LAYER M2 ;
        RECT 0.7 7.84 1.02 8.12 ;
  LAYER M2 ;
        RECT 1.55 17.92 2.75 18.2 ;
  LAYER M2 ;
        RECT 1.55 27.16 2.75 27.44 ;
  LAYER M2 ;
        RECT 1.56 17.92 1.88 18.2 ;
  LAYER M1 ;
        RECT 1.595 18.06 1.845 27.3 ;
  LAYER M2 ;
        RECT 1.56 27.16 1.88 27.44 ;
  LAYER M2 ;
        RECT 1.13 7.84 1.45 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.98 1.43 18.06 ;
  LAYER M2 ;
        RECT 1.29 17.92 1.72 18.2 ;
  LAYER M2 ;
        RECT 1.13 7.84 1.45 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.82 1.43 8.14 ;
  LAYER M2 ;
        RECT 1.13 17.92 1.45 18.2 ;
  LAYER M3 ;
        RECT 1.15 17.9 1.43 18.22 ;
  LAYER M2 ;
        RECT 1.13 7.84 1.45 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.82 1.43 8.14 ;
  LAYER M2 ;
        RECT 1.13 17.92 1.45 18.2 ;
  LAYER M3 ;
        RECT 1.15 17.9 1.43 18.22 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 1.29 2.8 2.58 3.08 ;
  LAYER M1 ;
        RECT 2.455 2.94 2.705 7.14 ;
  LAYER M2 ;
        RECT 2.58 7 3.87 7.28 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 7.14 4.01 7.98 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M1 ;
        RECT 2.455 7.14 2.705 12.18 ;
  LAYER M2 ;
        RECT 1.29 12.04 2.58 12.32 ;
  LAYER M1 ;
        RECT 2.455 2.855 2.705 3.025 ;
  LAYER M2 ;
        RECT 2.41 2.8 2.75 3.08 ;
  LAYER M1 ;
        RECT 2.455 7.055 2.705 7.225 ;
  LAYER M2 ;
        RECT 2.41 7 2.75 7.28 ;
  LAYER M1 ;
        RECT 2.455 2.855 2.705 3.025 ;
  LAYER M2 ;
        RECT 2.41 2.8 2.75 3.08 ;
  LAYER M1 ;
        RECT 2.455 7.055 2.705 7.225 ;
  LAYER M2 ;
        RECT 2.41 7 2.75 7.28 ;
  LAYER M1 ;
        RECT 2.455 2.855 2.705 3.025 ;
  LAYER M2 ;
        RECT 2.41 2.8 2.75 3.08 ;
  LAYER M1 ;
        RECT 2.455 7.055 2.705 7.225 ;
  LAYER M2 ;
        RECT 2.41 7 2.75 7.28 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 2.455 2.855 2.705 3.025 ;
  LAYER M2 ;
        RECT 2.41 2.8 2.75 3.08 ;
  LAYER M1 ;
        RECT 2.455 7.055 2.705 7.225 ;
  LAYER M2 ;
        RECT 2.41 7 2.75 7.28 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 2.455 2.855 2.705 3.025 ;
  LAYER M2 ;
        RECT 2.41 2.8 2.75 3.08 ;
  LAYER M1 ;
        RECT 2.455 7.055 2.705 7.225 ;
  LAYER M2 ;
        RECT 2.41 7 2.75 7.28 ;
  LAYER M1 ;
        RECT 2.455 12.095 2.705 12.265 ;
  LAYER M2 ;
        RECT 2.41 12.04 2.75 12.32 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 2.455 2.855 2.705 3.025 ;
  LAYER M2 ;
        RECT 2.41 2.8 2.75 3.08 ;
  LAYER M1 ;
        RECT 2.455 7.055 2.705 7.225 ;
  LAYER M2 ;
        RECT 2.41 7 2.75 7.28 ;
  LAYER M1 ;
        RECT 2.455 12.095 2.705 12.265 ;
  LAYER M2 ;
        RECT 2.41 12.04 2.75 12.32 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 2.455 18.815 2.705 22.345 ;
  LAYER M1 ;
        RECT 2.455 17.555 2.705 18.565 ;
  LAYER M1 ;
        RECT 2.455 15.455 2.705 16.465 ;
  LAYER M1 ;
        RECT 2.025 18.815 2.275 22.345 ;
  LAYER M1 ;
        RECT 2.885 18.815 3.135 22.345 ;
  LAYER M2 ;
        RECT 1.98 15.82 3.18 16.1 ;
  LAYER M2 ;
        RECT 1.98 21.7 3.18 21.98 ;
  LAYER M2 ;
        RECT 1.55 22.12 2.75 22.4 ;
  LAYER M2 ;
        RECT 1.55 17.92 2.75 18.2 ;
  LAYER M3 ;
        RECT 2.87 15.8 3.15 22 ;
  LAYER M1 ;
        RECT 2.455 23.015 2.705 26.545 ;
  LAYER M1 ;
        RECT 2.455 26.795 2.705 27.805 ;
  LAYER M1 ;
        RECT 2.455 28.895 2.705 29.905 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 26.545 ;
  LAYER M1 ;
        RECT 2.885 23.015 3.135 26.545 ;
  LAYER M2 ;
        RECT 1.98 29.26 3.18 29.54 ;
  LAYER M2 ;
        RECT 1.98 23.38 3.18 23.66 ;
  LAYER M2 ;
        RECT 1.55 22.96 2.75 23.24 ;
  LAYER M2 ;
        RECT 1.55 27.16 2.75 27.44 ;
  LAYER M3 ;
        RECT 2.87 23.36 3.15 29.56 ;
  END 
END MY_RO
