* SPICE3 file created from MY_OPAMP_0.ext - technology: sky130A

.subckt MY_OPAMP_0 Y VP VN A B
X0 li_1093_1495# m1_1258_1568# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.814e+12p ps=2.368e+07u w=2.1e+06u l=150000u
X1 VP m1_1258_1568# li_1093_1495# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X2 m1_1258_1568# m1_1258_1568# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X3 VP m1_1258_1568# m1_1258_1568# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X4 m1_516_1316# m1_1258_1568# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X5 VP m1_1258_1568# m1_516_1316# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X6 m1_946_1400# PMOS_4T_31631261_X1_Y1_1678560933_0/a_200_252# m1_516_1316# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X7 m1_516_1316# PMOS_4T_31631261_X1_Y1_1678560933_0/a_200_252# m1_946_1400# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X8 m1_570_1400# PMOS_4T_31631261_X1_Y1_1678560933_1/a_200_252# m1_516_1316# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X9 m1_516_1316# PMOS_4T_31631261_X1_Y1_1678560933_1/a_200_252# m1_570_1400# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X10 m1_946_1400# m1_570_1400# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X11 SUB m1_570_1400# m1_946_1400# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X12 m1_570_1400# m1_570_1400# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X13 SUB m1_570_1400# m1_570_1400# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X14 li_1093_1495# m1_946_1400# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X15 SUB m1_946_1400# li_1093_1495# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X16 m1_1258_1568# VP SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X17 SUB VP m1_1258_1568# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 Y m1_516_1316# 0.01fF
C1 m1_946_1400# m1_516_1316# 0.71fF
C2 B m1_516_1316# 0.01fF
C3 A m1_516_1316# 0.02fF
C4 li_1093_1495# m1_516_1316# 0.01fF
C5 PMOS_4T_31631261_X1_Y1_1678560933_0/a_200_252# VP 0.19fF
C6 VP m1_516_1316# 1.49fF
C7 m1_1258_1568# VN 0.02fF
C8 m1_570_1400# m1_516_1316# 0.87fF
C9 Y VN 0.08fF
C10 m1_946_1400# VN 0.21fF
C11 B VN 0.01fF
C12 A VN 0.00fF
C13 PMOS_4T_31631261_X1_Y1_1678560933_1/a_200_252# VP 0.19fF
C14 PMOS_4T_31631261_X1_Y1_1678560933_1/a_200_252# m1_570_1400# 0.04fF
C15 VP VN 0.34fF
C16 m1_1258_1568# Y 0.06fF
C17 m1_946_1400# m1_1258_1568# 0.29fF
C18 m1_570_1400# VN 0.06fF
C19 m1_1258_1568# B 0.01fF
C20 m1_946_1400# Y 0.08fF
C21 m1_1258_1568# A 0.02fF
C22 PMOS_4T_31631261_X1_Y1_1678560933_0/a_200_252# m1_516_1316# 0.03fF
C23 m1_1258_1568# li_1093_1495# 0.26fF
C24 Y B 0.00fF
C25 m1_946_1400# A 0.00fF
C26 m1_1258_1568# VP 2.92fF
C27 m1_946_1400# li_1093_1495# 0.14fF
C28 A B 0.04fF
C29 m1_570_1400# m1_1258_1568# 0.28fF
C30 VP Y 0.13fF
C31 m1_946_1400# VP 0.82fF
C32 m1_570_1400# Y 0.06fF
C33 m1_946_1400# m1_570_1400# 0.50fF
C34 VP B 0.05fF
C35 A VP 0.05fF
C36 PMOS_4T_31631261_X1_Y1_1678560933_1/a_200_252# m1_516_1316# 0.03fF
C37 m1_570_1400# B 0.07fF
C38 li_1093_1495# VP 0.73fF
C39 m1_570_1400# A 0.01fF
C40 m1_570_1400# li_1093_1495# 0.00fF
C41 VN m1_516_1316# 0.06fF
C42 m1_570_1400# VP 0.62fF
C43 m1_1258_1568# m1_516_1316# 0.23fF
C44 m1_946_1400# PMOS_4T_31631261_X1_Y1_1678560933_0/a_200_252# 0.04fF
C45 VP SUB 12.80fF
C46 li_1093_1495# SUB 1.15fF **FLOATING
C47 m1_570_1400# SUB 1.64fF **FLOATING
C48 PMOS_4T_31631261_X1_Y1_1678560933_1/a_200_252# SUB 0.25fF **FLOATING
C49 m1_946_1400# SUB 1.50fF **FLOATING
C50 m1_516_1316# SUB 0.22fF **FLOATING
C51 PMOS_4T_31631261_X1_Y1_1678560933_0/a_200_252# SUB 0.25fF **FLOATING
C52 m1_1258_1568# SUB 0.85fF **FLOATING
.ends
