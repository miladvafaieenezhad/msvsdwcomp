MACRO MY_FUNCTION
  ORIGIN 0 0 ;
  FOREIGN MY_FUNCTION 0 0 ;
  SIZE 15.48 BY 15.12 ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
      LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
      LAYER M2 ;
        RECT 9.3 2.8 9.62 3.08 ;
      LAYER M3 ;
        RECT 9.32 2.94 9.6 12.18 ;
      LAYER M2 ;
        RECT 9.3 12.04 9.62 12.32 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.72 2.38 10.92 2.66 ;
      LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
      LAYER M2 ;
        RECT 3.01 2.38 9.89 2.66 ;
      LAYER M1 ;
        RECT 2.885 2.52 3.135 12.18 ;
      LAYER M2 ;
        RECT 1.29 12.04 3.01 12.32 ;
    END
  END B
  PIN VP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 7.14 0.7 8.34 0.98 ;
      LAYER M2 ;
        RECT 12.3 0.7 13.5 0.98 ;
      LAYER M3 ;
        RECT 11.04 0.68 11.32 6.46 ;
      LAYER M2 ;
        RECT 13.16 14.14 14.36 14.42 ;
      LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
      LAYER M2 ;
        RECT 8.17 0.7 9.03 0.98 ;
      LAYER M1 ;
        RECT 8.905 0.84 9.155 1.26 ;
      LAYER M2 ;
        RECT 9.03 1.12 12.04 1.4 ;
      LAYER M1 ;
        RECT 11.915 0.84 12.165 1.26 ;
      LAYER M2 ;
        RECT 12.04 0.7 12.47 0.98 ;
      LAYER M2 ;
        RECT 11.02 1.12 11.34 1.4 ;
      LAYER M3 ;
        RECT 11.04 1.075 11.32 1.445 ;
      LAYER M3 ;
        RECT 11.04 6.3 11.32 13.86 ;
      LAYER M2 ;
        RECT 11.18 13.72 12.47 14 ;
      LAYER M1 ;
        RECT 12.345 13.86 12.595 14.28 ;
      LAYER M2 ;
        RECT 12.47 14.14 13.33 14.42 ;
      LAYER M2 ;
        RECT 8.17 13.72 11.18 14 ;
      LAYER M1 ;
        RECT 8.045 13.86 8.295 14.28 ;
      LAYER M2 ;
        RECT 7.31 14.14 8.17 14.42 ;
    END
  END VP
  PIN VN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M2 ;
        RECT 4.56 0.7 5.76 0.98 ;
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M2 ;
        RECT 8.86 14.14 10.06 14.42 ;
      LAYER M2 ;
        RECT 10.58 14.14 11.78 14.42 ;
      LAYER M3 ;
        RECT 1.58 1.075 1.86 1.445 ;
      LAYER M2 ;
        RECT 1.72 1.12 4.73 1.4 ;
      LAYER M3 ;
        RECT 4.59 0.84 4.87 1.26 ;
      LAYER M2 ;
        RECT 4.57 0.7 4.89 0.98 ;
      LAYER M3 ;
        RECT 1.58 6.72 1.86 8.4 ;
      LAYER M3 ;
        RECT 1.58 9.055 1.86 9.425 ;
      LAYER M2 ;
        RECT 1.72 9.1 3.44 9.38 ;
      LAYER M3 ;
        RECT 3.3 9.055 3.58 9.425 ;
      LAYER M3 ;
        RECT 3.3 13.675 3.58 14.045 ;
      LAYER M4 ;
        RECT 3.44 13.46 9.03 14.26 ;
      LAYER M3 ;
        RECT 8.89 13.86 9.17 14.28 ;
      LAYER M2 ;
        RECT 8.87 14.14 9.19 14.42 ;
      LAYER M2 ;
        RECT 9.89 14.14 10.75 14.42 ;
    END
  END VN
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
      LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
      LAYER M2 ;
        RECT 4.73 12.04 6.45 12.32 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.98 2.8 3.18 3.08 ;
      LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
      LAYER M2 ;
        RECT 3.01 2.8 3.87 3.08 ;
      LAYER M1 ;
        RECT 3.745 2.94 3.995 3.36 ;
      LAYER M2 ;
        RECT 3.87 3.22 10.75 3.5 ;
      LAYER M3 ;
        RECT 10.61 2.94 10.89 3.36 ;
      LAYER M2 ;
        RECT 10.75 2.8 12.47 3.08 ;
    END
  END F
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
      LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
      LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
      LAYER M2 ;
        RECT 10.58 7.84 11.78 8.12 ;
      LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
      LAYER M2 ;
        RECT 5.59 7 7.31 7.28 ;
      LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
      LAYER M3 ;
        RECT 8.03 7.14 8.31 7.98 ;
      LAYER M2 ;
        RECT 8.17 7.84 9.03 8.12 ;
      LAYER M2 ;
        RECT 9.89 7.84 10.75 8.12 ;
      LAYER M2 ;
        RECT 11.61 7.84 12.47 8.12 ;
      LAYER M1 ;
        RECT 12.345 7.14 12.595 7.98 ;
      LAYER M2 ;
        RECT 12.31 7 12.63 7.28 ;
    END
  END Y
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 10.58 12.04 11.78 12.32 ;
      LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
      LAYER M2 ;
        RECT 11.61 12.04 13.33 12.32 ;
    END
  END C
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 4.56 2.8 5.76 3.08 ;
      LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
      LAYER M2 ;
        RECT 5.59 2.8 7.31 3.08 ;
    END
  END E
  OBS 
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 13.59 8.26 14.79 8.54 ;
  LAYER M2 ;
        RECT 9.89 7 11.61 7.28 ;
  LAYER M1 ;
        RECT 11.485 7.14 11.735 7.56 ;
  LAYER M2 ;
        RECT 11.61 7.42 12.9 7.7 ;
  LAYER M1 ;
        RECT 12.775 7.56 13.025 8.4 ;
  LAYER M2 ;
        RECT 12.9 8.26 13.76 8.54 ;
  LAYER M1 ;
        RECT 11.485 7.055 11.735 7.225 ;
  LAYER M2 ;
        RECT 11.44 7 11.78 7.28 ;
  LAYER M1 ;
        RECT 11.485 7.475 11.735 7.645 ;
  LAYER M2 ;
        RECT 11.44 7.42 11.78 7.7 ;
  LAYER M1 ;
        RECT 12.775 7.475 13.025 7.645 ;
  LAYER M2 ;
        RECT 12.73 7.42 13.07 7.7 ;
  LAYER M1 ;
        RECT 12.775 8.315 13.025 8.485 ;
  LAYER M2 ;
        RECT 12.73 8.26 13.07 8.54 ;
  LAYER M1 ;
        RECT 11.485 7.055 11.735 7.225 ;
  LAYER M2 ;
        RECT 11.44 7 11.78 7.28 ;
  LAYER M1 ;
        RECT 11.485 7.475 11.735 7.645 ;
  LAYER M2 ;
        RECT 11.44 7.42 11.78 7.7 ;
  LAYER M1 ;
        RECT 12.775 7.475 13.025 7.645 ;
  LAYER M2 ;
        RECT 12.73 7.42 13.07 7.7 ;
  LAYER M1 ;
        RECT 12.775 8.315 13.025 8.485 ;
  LAYER M2 ;
        RECT 12.73 8.26 13.07 8.54 ;
  LAYER M2 ;
        RECT 9.72 6.58 10.92 6.86 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 8.6 6.58 9.89 6.86 ;
  LAYER M1 ;
        RECT 8.475 6.72 8.725 7.56 ;
  LAYER M2 ;
        RECT 7.31 7.42 8.6 7.7 ;
  LAYER M1 ;
        RECT 7.185 7.56 7.435 8.4 ;
  LAYER M2 ;
        RECT 6.88 8.26 7.31 8.54 ;
  LAYER M1 ;
        RECT 7.185 7.475 7.435 7.645 ;
  LAYER M2 ;
        RECT 7.14 7.42 7.48 7.7 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 8.485 ;
  LAYER M2 ;
        RECT 7.14 8.26 7.48 8.54 ;
  LAYER M1 ;
        RECT 8.475 6.635 8.725 6.805 ;
  LAYER M2 ;
        RECT 8.43 6.58 8.77 6.86 ;
  LAYER M1 ;
        RECT 8.475 7.475 8.725 7.645 ;
  LAYER M2 ;
        RECT 8.43 7.42 8.77 7.7 ;
  LAYER M1 ;
        RECT 7.185 7.475 7.435 7.645 ;
  LAYER M2 ;
        RECT 7.14 7.42 7.48 7.7 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 8.485 ;
  LAYER M2 ;
        RECT 7.14 8.26 7.48 8.54 ;
  LAYER M1 ;
        RECT 8.475 6.635 8.725 6.805 ;
  LAYER M2 ;
        RECT 8.43 6.58 8.77 6.86 ;
  LAYER M1 ;
        RECT 8.475 7.475 8.725 7.645 ;
  LAYER M2 ;
        RECT 8.43 7.42 8.77 7.7 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M2 ;
        RECT 1.29 7.84 3.87 8.12 ;
  LAYER M2 ;
        RECT 4.73 7.84 5.59 8.12 ;
  LAYER M1 ;
        RECT 5.465 7.98 5.715 8.82 ;
  LAYER M2 ;
        RECT 5.59 8.68 8.17 8.96 ;
  LAYER M1 ;
        RECT 8.045 8.4 8.295 8.82 ;
  LAYER M2 ;
        RECT 8.17 8.26 8.6 8.54 ;
  LAYER M2 ;
        RECT 9.46 8.26 11.18 8.54 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.065 ;
  LAYER M2 ;
        RECT 5.42 7.84 5.76 8.12 ;
  LAYER M1 ;
        RECT 5.465 8.735 5.715 8.905 ;
  LAYER M2 ;
        RECT 5.42 8.68 5.76 8.96 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 8.485 ;
  LAYER M2 ;
        RECT 8 8.26 8.34 8.54 ;
  LAYER M1 ;
        RECT 8.045 8.735 8.295 8.905 ;
  LAYER M2 ;
        RECT 8 8.68 8.34 8.96 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.065 ;
  LAYER M2 ;
        RECT 5.42 7.84 5.76 8.12 ;
  LAYER M1 ;
        RECT 5.465 8.735 5.715 8.905 ;
  LAYER M2 ;
        RECT 5.42 8.68 5.76 8.96 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 8.485 ;
  LAYER M2 ;
        RECT 8 8.26 8.34 8.54 ;
  LAYER M1 ;
        RECT 8.045 8.735 8.295 8.905 ;
  LAYER M2 ;
        RECT 8 8.68 8.34 8.96 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.065 ;
  LAYER M2 ;
        RECT 5.42 7.84 5.76 8.12 ;
  LAYER M1 ;
        RECT 5.465 8.735 5.715 8.905 ;
  LAYER M2 ;
        RECT 5.42 8.68 5.76 8.96 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 8.485 ;
  LAYER M2 ;
        RECT 8 8.26 8.34 8.54 ;
  LAYER M1 ;
        RECT 8.045 8.735 8.295 8.905 ;
  LAYER M2 ;
        RECT 8 8.68 8.34 8.96 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.065 ;
  LAYER M2 ;
        RECT 5.42 7.84 5.76 8.12 ;
  LAYER M1 ;
        RECT 5.465 8.735 5.715 8.905 ;
  LAYER M2 ;
        RECT 5.42 8.68 5.76 8.96 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 8.485 ;
  LAYER M2 ;
        RECT 8 8.26 8.34 8.54 ;
  LAYER M1 ;
        RECT 8.045 8.735 8.295 8.905 ;
  LAYER M2 ;
        RECT 8 8.68 8.34 8.96 ;
  LAYER M2 ;
        RECT 1.98 7 3.18 7.28 ;
  LAYER M2 ;
        RECT 4.13 6.58 5.33 6.86 ;
  LAYER M2 ;
        RECT 3.01 7 3.87 7.28 ;
  LAYER M1 ;
        RECT 3.745 6.72 3.995 7.14 ;
  LAYER M2 ;
        RECT 3.87 6.58 4.3 6.86 ;
  LAYER M1 ;
        RECT 3.745 6.635 3.995 6.805 ;
  LAYER M2 ;
        RECT 3.7 6.58 4.04 6.86 ;
  LAYER M1 ;
        RECT 3.745 7.055 3.995 7.225 ;
  LAYER M2 ;
        RECT 3.7 7 4.04 7.28 ;
  LAYER M1 ;
        RECT 3.745 6.635 3.995 6.805 ;
  LAYER M2 ;
        RECT 3.7 6.58 4.04 6.86 ;
  LAYER M1 ;
        RECT 3.745 7.055 3.995 7.225 ;
  LAYER M2 ;
        RECT 3.7 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 12.73 6.58 13.93 6.86 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.72 7.45 7.98 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.3 7.88 6.72 ;
  LAYER M4 ;
        RECT 7.74 5.9 11.61 6.7 ;
  LAYER M3 ;
        RECT 11.47 6.3 11.75 6.72 ;
  LAYER M2 ;
        RECT 11.61 6.58 12.9 6.86 ;
  LAYER M2 ;
        RECT 13.17 6.58 13.49 6.86 ;
  LAYER M3 ;
        RECT 13.19 6.72 13.47 7.98 ;
  LAYER M2 ;
        RECT 13.17 7.84 13.49 8.12 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.56 11.75 6.88 ;
  LAYER M3 ;
        RECT 7.6 6.115 7.88 6.485 ;
  LAYER M4 ;
        RECT 7.575 5.9 7.905 6.7 ;
  LAYER M3 ;
        RECT 11.47 6.115 11.75 6.485 ;
  LAYER M4 ;
        RECT 11.445 5.9 11.775 6.7 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.56 11.75 6.88 ;
  LAYER M3 ;
        RECT 7.6 6.115 7.88 6.485 ;
  LAYER M4 ;
        RECT 7.575 5.9 7.905 6.7 ;
  LAYER M3 ;
        RECT 11.47 6.115 11.75 6.485 ;
  LAYER M4 ;
        RECT 11.445 5.9 11.775 6.7 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.56 11.75 6.88 ;
  LAYER M2 ;
        RECT 13.17 6.58 13.49 6.86 ;
  LAYER M3 ;
        RECT 13.19 6.56 13.47 6.88 ;
  LAYER M2 ;
        RECT 13.17 7.84 13.49 8.12 ;
  LAYER M3 ;
        RECT 13.19 7.82 13.47 8.14 ;
  LAYER M3 ;
        RECT 7.6 6.115 7.88 6.485 ;
  LAYER M4 ;
        RECT 7.575 5.9 7.905 6.7 ;
  LAYER M3 ;
        RECT 11.47 6.115 11.75 6.485 ;
  LAYER M4 ;
        RECT 11.445 5.9 11.775 6.7 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.56 11.75 6.88 ;
  LAYER M2 ;
        RECT 13.17 6.58 13.49 6.86 ;
  LAYER M3 ;
        RECT 13.19 6.56 13.47 6.88 ;
  LAYER M2 ;
        RECT 13.17 7.84 13.49 8.12 ;
  LAYER M3 ;
        RECT 13.19 7.82 13.47 8.14 ;
  LAYER M3 ;
        RECT 7.6 6.115 7.88 6.485 ;
  LAYER M4 ;
        RECT 7.575 5.9 7.905 6.7 ;
  LAYER M3 ;
        RECT 11.47 6.115 11.75 6.485 ;
  LAYER M4 ;
        RECT 11.445 5.9 11.775 6.7 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 9.72 0.7 11.35 0.98 ;
  LAYER M2 ;
        RECT 9.29 6.16 11.35 6.44 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 9.72 6.58 10.92 6.86 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M2 ;
        RECT 9.72 2.38 10.92 2.66 ;
  LAYER M3 ;
        RECT 11.04 0.68 11.32 6.46 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 1.55 0.7 2.75 0.98 ;
  LAYER M2 ;
        RECT 1.55 6.58 2.75 6.86 ;
  LAYER M2 ;
        RECT 1.98 7 3.18 7.28 ;
  LAYER M2 ;
        RECT 1.98 2.8 3.18 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M2 ;
        RECT 8.86 14.14 10.06 14.42 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M2 ;
        RECT 10.58 14.14 11.78 14.42 ;
  LAYER M2 ;
        RECT 10.58 7.84 11.78 8.12 ;
  LAYER M2 ;
        RECT 10.58 12.04 11.78 12.32 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 4.56 0.7 5.76 0.98 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 4.56 2.8 5.76 3.08 ;
  LAYER M2 ;
        RECT 4.13 6.58 5.33 6.86 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 7.14 0.7 8.34 0.98 ;
  LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M2 ;
        RECT 12.3 0.7 13.5 0.98 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
  LAYER M2 ;
        RECT 12.73 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M2 ;
        RECT 13.16 14.14 14.36 14.42 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
  LAYER M2 ;
        RECT 13.59 8.26 14.79 8.54 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  END 
END MY_FUNCTION
