* SPICE3 file created from MY_RO_0.ext - technology: sky130A

.subckt MY_RO_0 VN VP A Y
X0 INV_51706272_0_0_1677482275_0/m1_312_1400# m1_226_1568# m1_312_4508# m1_312_4508# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 m1_312_4508# m1_226_1568# INV_51706272_0_0_1677482275_0/m1_312_1400# m1_312_4508# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 INV_51706272_0_0_1677482275_0/m1_312_1400# m1_226_1568# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 SUB m1_226_1568# INV_51706272_0_0_1677482275_0/m1_312_1400# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 m1_226_1568# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# m1_312_4508# m1_312_4508# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 m1_312_4508# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# m1_226_1568# m1_312_4508# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# m1_312_4508# m1_312_4508# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 m1_312_4508# STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# m1_312_4508# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 SUB STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 m1_226_1568# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 SUB STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# m1_226_1568# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# 0.35fF
C1 INV_51706272_0_0_1677482275_0/m1_312_1400# m1_226_1568# 0.13fF
C2 Y STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# 0.00fF
C3 A m1_226_1568# 0.00fF
C4 INV_51706272_0_0_1677482275_0/m1_312_1400# m1_312_4508# 0.70fF
C5 m1_226_1568# VP 0.92fF
C6 STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# m1_226_1568# 0.01fF
C7 VP m1_312_4508# 0.00fF
C8 m1_226_1568# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# 0.18fF
C9 STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# m1_312_4508# 0.55fF
C10 m1_312_4508# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# 1.57fF
C11 Y m1_312_4508# 0.40fF
C12 A VN 0.01fF
C13 INV_51706272_0_0_1677482275_0/m1_312_1400# VP 0.00fF
C14 VP VN 0.94fF
C15 m1_226_1568# m1_312_4508# 1.72fF
C16 INV_51706272_0_0_1677482275_0/m1_312_1400# STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# 0.00fF
C17 VN STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# 0.26fF
C18 Y VP 0.00fF
C19 VP SUB 0.28fF
C20 STAGE2_INV_5734008_0_0_1677482276_0/m1_828_560# SUB 1.45fF **FLOATING
C21 m1_226_1568# SUB 2.98fF **FLOATING
C22 STAGE2_INV_5734008_0_0_1677482276_0/li_491_571# SUB 2.37fF **FLOATING
C23 m1_312_4508# SUB 9.43fF **FLOATING
C24 INV_51706272_0_0_1677482275_0/m1_312_1400# SUB 0.80fF **FLOATING
.ends
