magic
tech sky130A
timestamp 1675936227
<< nwell >>
rect -210 -25 -5 165
<< nmos >>
rect -90 -215 -75 -65
<< pmos >>
rect -90 -5 -75 145
<< ndiff >>
rect -140 -80 -90 -65
rect -140 -200 -125 -80
rect -105 -200 -90 -80
rect -140 -215 -90 -200
rect -75 -80 -25 -65
rect -75 -200 -60 -80
rect -40 -200 -25 -80
rect -75 -215 -25 -200
<< pdiff >>
rect -140 130 -90 145
rect -140 10 -125 130
rect -105 10 -90 130
rect -140 -5 -90 10
rect -75 130 -25 145
rect -75 10 -60 130
rect -40 10 -25 130
rect -75 -5 -25 10
<< ndiffc >>
rect -125 -200 -105 -80
rect -60 -200 -40 -80
<< pdiffc >>
rect -125 10 -105 130
rect -60 10 -40 130
<< psubdiff >>
rect -190 -80 -140 -65
rect -190 -200 -175 -80
rect -155 -200 -140 -80
rect -190 -215 -140 -200
<< nsubdiff >>
rect -190 130 -140 145
rect -190 10 -175 130
rect -155 10 -140 130
rect -190 -5 -140 10
<< psubdiffcont >>
rect -175 -200 -155 -80
<< nsubdiffcont >>
rect -175 10 -155 130
<< poly >>
rect -90 145 -75 160
rect -90 -65 -75 -5
rect -90 -230 -75 -215
rect -115 -240 -75 -230
rect -115 -260 -105 -240
rect -85 -260 -75 -240
rect -115 -270 -75 -260
<< polycont >>
rect -105 -260 -85 -240
<< locali >>
rect -180 130 -95 140
rect -180 10 -175 130
rect -155 10 -125 130
rect -105 10 -95 130
rect -180 0 -95 10
rect -70 130 -30 140
rect -70 10 -60 130
rect -40 10 -30 130
rect -70 0 -30 10
rect -50 -70 -30 0
rect -180 -80 -95 -70
rect -180 -200 -175 -80
rect -155 -200 -125 -80
rect -105 -200 -95 -80
rect -180 -210 -95 -200
rect -70 -80 -30 -70
rect -70 -200 -60 -80
rect -40 -200 -30 -80
rect -70 -210 -30 -200
rect -50 -230 -30 -210
rect -210 -240 -75 -230
rect -210 -250 -105 -240
rect -115 -260 -105 -250
rect -85 -260 -75 -240
rect -50 -250 -5 -230
rect -115 -270 -75 -260
<< viali >>
rect -175 10 -155 130
rect -125 10 -105 130
rect -175 -200 -155 -80
rect -125 -200 -105 -80
<< metal1 >>
rect -210 130 -5 140
rect -210 10 -175 130
rect -155 10 -125 130
rect -105 10 -5 130
rect -210 0 -5 10
rect -210 -80 -5 -70
rect -210 -200 -175 -80
rect -155 -200 -125 -80
rect -105 -200 -5 -80
rect -210 -210 -5 -200
<< labels >>
rlabel locali -5 -240 -5 -240 3 Y
port 2 e
rlabel locali -210 -240 -210 -240 7 A
port 1 w
rlabel metal1 -210 75 -210 75 7 VP
port 3 w
rlabel metal1 -210 -140 -210 -140 7 VN
port 4 w
<< end >>
