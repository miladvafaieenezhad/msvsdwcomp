* SPICE3 file created from MY_INVERTER_0.ext - technology: sky130A

.subckt MY_INVERTER_0 A VN VP Y
X0 INV_72761973_0_0_1676281181_0/m1_312_1400# INV_72761973_0_0_1676281181_0/li_405_571# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 SUB INV_72761973_0_0_1676281181_0/li_405_571# INV_72761973_0_0_1676281181_0/m1_312_1400# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 INV_72761973_0_0_1676281181_0/m1_312_1400# INV_72761973_0_0_1676281181_0/li_405_571# INV_72761973_0_0_1676281181_0/PMOS_S_99486525_X1_Y1_1676281182_1676281181_0/w_0_0# INV_72761973_0_0_1676281181_0/PMOS_S_99486525_X1_Y1_1676281182_1676281181_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 INV_72761973_0_0_1676281181_0/PMOS_S_99486525_X1_Y1_1676281182_1676281181_0/w_0_0# INV_72761973_0_0_1676281181_0/li_405_571# INV_72761973_0_0_1676281181_0/m1_312_1400# INV_72761973_0_0_1676281181_0/PMOS_S_99486525_X1_Y1_1676281182_1676281181_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 INV_72761973_0_0_1676281181_0/PMOS_S_99486525_X1_Y1_1676281182_1676281181_0/w_0_0# SUB 3.18fF **FLOATING
.ends
