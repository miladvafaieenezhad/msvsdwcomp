MACRO MY_OPAMP
  ORIGIN 0 0 ;
  FOREIGN MY_OPAMP 0 0 ;
  SIZE 9.46 BY 15.12 ;
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 4.56 7.84 5.76 8.12 ;
      LAYER M2 ;
        RECT 7.14 8.26 8.34 8.54 ;
      LAYER M2 ;
        RECT 5.43 7.84 5.75 8.12 ;
      LAYER M1 ;
        RECT 5.465 7.56 5.715 7.98 ;
      LAYER M2 ;
        RECT 5.59 7.42 6.45 7.7 ;
      LAYER M1 ;
        RECT 6.325 7.56 6.575 8.4 ;
      LAYER M2 ;
        RECT 6.45 8.26 7.31 8.54 ;
    END
  END Y
  PIN VP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.98 0.7 3.18 0.98 ;
      LAYER M2 ;
        RECT 3.7 0.7 4.9 0.98 ;
      LAYER M3 ;
        RECT 1.15 8.66 1.43 14.44 ;
      LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
      LAYER M3 ;
        RECT 1.15 11.155 1.43 11.525 ;
      LAYER M2 ;
        RECT 1.29 11.2 4.3 11.48 ;
      LAYER M3 ;
        RECT 4.16 11.155 4.44 11.525 ;
      LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
      LAYER M2 ;
        RECT 3.01 0.7 3.87 0.98 ;
      LAYER M2 ;
        RECT 4.14 0.7 4.46 0.98 ;
      LAYER M3 ;
        RECT 4.16 0.84 4.44 8.4 ;
      LAYER M3 ;
        RECT 4.16 12.415 4.44 12.785 ;
      LAYER M2 ;
        RECT 4.3 12.46 6.45 12.74 ;
      LAYER M1 ;
        RECT 6.325 12.18 6.575 12.6 ;
      LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
    END
  END VP
  PIN VN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 8.03 0.68 8.31 6.46 ;
      LAYER M3 ;
        RECT 8.46 8.66 8.74 14.44 ;
      LAYER M3 ;
        RECT 8.03 6.3 8.31 7.56 ;
      LAYER M2 ;
        RECT 8.17 7.42 8.6 7.7 ;
      LAYER M3 ;
        RECT 8.46 7.56 8.74 8.82 ;
    END
  END VN
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.98 2.8 3.18 3.08 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
    END
  END B
  OBS 
  LAYER M3 ;
        RECT 2.01 7.82 2.29 12.34 ;
  LAYER M2 ;
        RECT 4.56 12.04 5.76 12.32 ;
  LAYER M3 ;
        RECT 2.01 11.575 2.29 11.945 ;
  LAYER M2 ;
        RECT 2.15 11.62 3.87 11.9 ;
  LAYER M1 ;
        RECT 3.745 11.76 3.995 12.18 ;
  LAYER M2 ;
        RECT 3.87 12.04 4.73 12.32 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M3 ;
        RECT 2.01 8.635 2.29 9.005 ;
  LAYER M4 ;
        RECT 2.15 8.42 6.45 9.22 ;
  LAYER M3 ;
        RECT 6.31 7.98 6.59 8.82 ;
  LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
  LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
  LAYER M3 ;
        RECT 6.31 7.82 6.59 8.14 ;
  LAYER M3 ;
        RECT 2.01 8.635 2.29 9.005 ;
  LAYER M4 ;
        RECT 1.985 8.42 2.315 9.22 ;
  LAYER M3 ;
        RECT 6.31 8.635 6.59 9.005 ;
  LAYER M4 ;
        RECT 6.285 8.42 6.615 9.22 ;
  LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
  LAYER M3 ;
        RECT 6.31 7.82 6.59 8.14 ;
  LAYER M3 ;
        RECT 2.01 8.635 2.29 9.005 ;
  LAYER M4 ;
        RECT 1.985 8.42 2.315 9.22 ;
  LAYER M3 ;
        RECT 6.31 8.635 6.59 9.005 ;
  LAYER M4 ;
        RECT 6.285 8.42 6.615 9.22 ;
  LAYER M2 ;
        RECT 1.55 6.58 2.75 6.86 ;
  LAYER M2 ;
        RECT 1.12 8.26 2.32 8.54 ;
  LAYER M2 ;
        RECT 4.13 6.58 5.33 6.86 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.72 1.86 8.4 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M2 ;
        RECT 2.58 6.58 4.3 6.86 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.98 7 3.18 7.28 ;
  LAYER M3 ;
        RECT 7.17 2.78 7.45 7.3 ;
  LAYER M2 ;
        RECT 2.85 7 3.17 7.28 ;
  LAYER M3 ;
        RECT 2.87 6.3 3.15 7.14 ;
  LAYER M4 ;
        RECT 3.01 5.9 7.31 6.7 ;
  LAYER M3 ;
        RECT 7.17 6.115 7.45 6.485 ;
  LAYER M2 ;
        RECT 2.85 7 3.17 7.28 ;
  LAYER M3 ;
        RECT 2.87 6.98 3.15 7.3 ;
  LAYER M3 ;
        RECT 2.87 6.115 3.15 6.485 ;
  LAYER M4 ;
        RECT 2.845 5.9 3.175 6.7 ;
  LAYER M3 ;
        RECT 7.17 6.115 7.45 6.485 ;
  LAYER M4 ;
        RECT 7.145 5.9 7.475 6.7 ;
  LAYER M2 ;
        RECT 2.85 7 3.17 7.28 ;
  LAYER M3 ;
        RECT 2.87 6.98 3.15 7.3 ;
  LAYER M3 ;
        RECT 2.87 6.115 3.15 6.485 ;
  LAYER M4 ;
        RECT 2.845 5.9 3.175 6.7 ;
  LAYER M3 ;
        RECT 7.17 6.115 7.45 6.485 ;
  LAYER M4 ;
        RECT 7.145 5.9 7.475 6.7 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 7.14 6.58 8.34 6.86 ;
  LAYER M2 ;
        RECT 7.14 12.46 8.34 12.74 ;
  LAYER M2 ;
        RECT 4.73 7 5.59 7.28 ;
  LAYER M3 ;
        RECT 5.45 7.14 5.73 7.56 ;
  LAYER M4 ;
        RECT 5.59 7.16 6.88 7.96 ;
  LAYER M3 ;
        RECT 6.74 6.72 7.02 7.56 ;
  LAYER M2 ;
        RECT 6.88 6.58 7.31 6.86 ;
  LAYER M3 ;
        RECT 6.74 7.56 7.02 11.76 ;
  LAYER M2 ;
        RECT 6.88 11.62 7.31 11.9 ;
  LAYER M3 ;
        RECT 7.17 11.76 7.45 12.6 ;
  LAYER M2 ;
        RECT 7.15 12.46 7.47 12.74 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 7.3 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M3 ;
        RECT 6.74 7.375 7.02 7.745 ;
  LAYER M4 ;
        RECT 6.715 7.16 7.045 7.96 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 7.3 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M3 ;
        RECT 6.74 7.375 7.02 7.745 ;
  LAYER M4 ;
        RECT 6.715 7.16 7.045 7.96 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 7.3 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M2 ;
        RECT 6.72 11.62 7.04 11.9 ;
  LAYER M3 ;
        RECT 6.74 11.6 7.02 11.92 ;
  LAYER M2 ;
        RECT 7.15 11.62 7.47 11.9 ;
  LAYER M3 ;
        RECT 7.17 11.6 7.45 11.92 ;
  LAYER M2 ;
        RECT 7.15 12.46 7.47 12.74 ;
  LAYER M3 ;
        RECT 7.17 12.44 7.45 12.76 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M3 ;
        RECT 6.74 7.375 7.02 7.745 ;
  LAYER M4 ;
        RECT 6.715 7.16 7.045 7.96 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 7.3 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M2 ;
        RECT 6.72 11.62 7.04 11.9 ;
  LAYER M3 ;
        RECT 6.74 11.6 7.02 11.92 ;
  LAYER M2 ;
        RECT 7.15 11.62 7.47 11.9 ;
  LAYER M3 ;
        RECT 7.17 11.6 7.45 11.92 ;
  LAYER M2 ;
        RECT 7.15 12.46 7.47 12.74 ;
  LAYER M3 ;
        RECT 7.17 12.44 7.45 12.76 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M3 ;
        RECT 6.74 7.375 7.02 7.745 ;
  LAYER M4 ;
        RECT 6.715 7.16 7.045 7.96 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 1.98 7.84 3.18 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 1.12 14.14 2.32 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.68 2.75 8.96 ;
  LAYER M3 ;
        RECT 2.01 7.82 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.12 8.26 2.32 8.54 ;
  LAYER M3 ;
        RECT 1.15 8.66 1.43 14.44 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 14.785 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 4.13 14.14 5.33 14.42 ;
  LAYER M2 ;
        RECT 4.13 8.26 5.33 8.54 ;
  LAYER M2 ;
        RECT 4.56 7.84 5.76 8.12 ;
  LAYER M2 ;
        RECT 4.56 12.04 5.76 12.32 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M2 ;
        RECT 7.14 0.7 8.34 0.98 ;
  LAYER M2 ;
        RECT 6.71 6.16 8.77 6.44 ;
  LAYER M3 ;
        RECT 7.17 2.78 7.45 7.3 ;
  LAYER M2 ;
        RECT 7.14 6.58 8.34 6.86 ;
  LAYER M3 ;
        RECT 8.03 0.68 8.31 6.46 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M2 ;
        RECT 7.14 14.14 8.77 14.42 ;
  LAYER M2 ;
        RECT 6.71 8.68 8.77 8.96 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 7.14 8.26 8.34 8.54 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 7.14 12.46 8.34 12.74 ;
  LAYER M3 ;
        RECT 8.46 8.66 8.74 14.44 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 1.98 0.7 3.18 0.98 ;
  LAYER M2 ;
        RECT 1.98 7 3.18 7.28 ;
  LAYER M2 ;
        RECT 1.98 2.8 3.18 3.08 ;
  LAYER M2 ;
        RECT 1.55 6.58 2.75 6.86 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M2 ;
        RECT 3.7 0.7 4.9 0.98 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 4.13 6.58 5.33 6.86 ;
  END 
END MY_OPAMP
