.subckt inverter  A VP Y VN
XM1 Y A VN VN sky130_fd_pr__nfet_01v8 w=14.7e-7 l=150e-9 nf=2 m=1
XM2 Y A VP VP sky130_fd_pr__pfet_01v8 w=14.7e-7 l=150e-9  nf=2 m=1
.ends inverter

