** sch_path: /home/milad/.xschem/xschem_library/VSD/week3/(3)post_layout_ring/RO_test.sch
**.subckt RO_test
Vdd VDD GND 1.8
x1 VA VDD VA GND 3_stages_RO
**** begin user architecture code


.include ~/.xschem/xschem_library/VSD/week3/(3)post_layout_ring/MY_RO.spice
.IC v(VA)=1.8
.tran 0.1n 15n
.measure tran T  TRIG v(Va) TD=5n VAL=0.9 FALL=1  TARG v(Va) TD=5n VAL=0.9 FALL=2
.save all

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
