* SPICE3 file created from MY_OPAMP_0.ext - technology: sky130A

.subckt MY_OPAMP_0 Y VP VN A B
X0 li_1093_1495# m1_946_1400# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 SUB m1_946_1400# li_1093_1495# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 m1_1258_1568# VP SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 SUB VP m1_1258_1568# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 li_1093_1495# m1_1258_1568# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.628e+11p ps=6.88e+06u w=420000u l=150000u
X5 VP m1_1258_1568# li_1093_1495# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VP m1_1258_1568# m1_516_1316# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 m1_1258_1568# m1_1258_1568# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VP m1_1258_1568# m1_1258_1568# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 m1_516_1316# m1_1258_1568# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 m1_946_1400# m1_570_1400# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 SUB m1_570_1400# m1_946_1400# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 m1_570_1400# m1_570_1400# SUB SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 SUB m1_570_1400# m1_570_1400# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 m1_946_1400# PMOS_4T_68898473_X1_Y1_1678026281_0/a_200_252# m1_516_1316# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 m1_516_1316# PMOS_4T_68898473_X1_Y1_1678026281_0/a_200_252# m1_946_1400# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 m1_570_1400# PMOS_4T_68898473_X1_Y1_1678026281_1/a_200_252# m1_516_1316# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 m1_516_1316# PMOS_4T_68898473_X1_Y1_1678026281_1/a_200_252# m1_570_1400# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 PMOS_4T_68898473_X1_Y1_1678026281_1/a_200_252# m1_516_1316# 0.03fF
C1 Y VN 0.08fF
C2 Y m1_1258_1568# 0.06fF
C3 Y VP 0.12fF
C4 Y m1_570_1400# 0.06fF
C5 m1_516_1316# B 0.01fF
C6 m1_516_1316# m1_946_1400# 0.67fF
C7 m1_1258_1568# li_1093_1495# 0.25fF
C8 VP li_1093_1495# 0.70fF
C9 li_1093_1495# m1_570_1400# 0.00fF
C10 m1_1258_1568# VN 0.02fF
C11 VP VN 0.34fF
C12 VN m1_570_1400# 0.06fF
C13 m1_1258_1568# VP 2.99fF
C14 m1_1258_1568# m1_570_1400# 0.27fF
C15 A VN 0.01fF
C16 VP PMOS_4T_68898473_X1_Y1_1678026281_0/a_200_252# 0.23fF
C17 A m1_1258_1568# 0.02fF
C18 VP m1_570_1400# 0.61fF
C19 A VP 0.06fF
C20 A m1_570_1400# 0.01fF
C21 Y B 0.00fF
C22 Y m1_946_1400# 0.07fF
C23 Y m1_516_1316# 0.00fF
C24 li_1093_1495# m1_946_1400# 0.14fF
C25 li_1093_1495# m1_516_1316# 0.01fF
C26 VP PMOS_4T_68898473_X1_Y1_1678026281_1/a_200_252# 0.23fF
C27 PMOS_4T_68898473_X1_Y1_1678026281_1/a_200_252# m1_570_1400# 0.04fF
C28 VN B 0.01fF
C29 m1_1258_1568# B 0.01fF
C30 VN m1_946_1400# 0.21fF
C31 m1_1258_1568# m1_946_1400# 0.29fF
C32 VP B 0.05fF
C33 m1_946_1400# PMOS_4T_68898473_X1_Y1_1678026281_0/a_200_252# 0.04fF
C34 B m1_570_1400# 0.08fF
C35 m1_516_1316# VN 0.07fF
C36 VP m1_946_1400# 0.86fF
C37 A B 0.06fF
C38 m1_946_1400# m1_570_1400# 0.49fF
C39 m1_1258_1568# m1_516_1316# 0.22fF
C40 A m1_946_1400# 0.00fF
C41 m1_516_1316# PMOS_4T_68898473_X1_Y1_1678026281_0/a_200_252# 0.03fF
C42 VP m1_516_1316# 1.50fF
C43 m1_516_1316# m1_570_1400# 0.81fF
C44 A m1_516_1316# 0.02fF
C45 VP SUB 12.92fF
C46 m1_570_1400# SUB 1.74fF **FLOATING
C47 PMOS_4T_68898473_X1_Y1_1678026281_1/a_200_252# SUB 0.42fF **FLOATING
C48 m1_946_1400# SUB 1.57fF **FLOATING
C49 m1_516_1316# SUB 0.26fF **FLOATING
C50 PMOS_4T_68898473_X1_Y1_1678026281_0/a_200_252# SUB 0.42fF **FLOATING
C51 m1_1258_1568# SUB 1.03fF **FLOATING
C52 li_1093_1495# SUB 1.15fF **FLOATING
.ends
